Simple MOS Current Mirror

.INCLUDE simple_mos_current_mirror_simulation_netlist.spice

* Interactive simulation main entry *
.CONTROL

* Make a directory for our output simulation files.
shell mkdir -p results 
* Generic prefix for our output files
set generic_prefix = 'results/simple_mos_current_mirror_simulation'

echo  '* Operating point analysis: Current match '

OP                      
print all               
* Output current over constant input current (with 1V load): should be 1 for best match.
print (v2#branch/v1#branch)

echo '* DC analysis: Voltage dependence of current mirror'

DC V2 0V 3V 0.1V          ; Sweep Drain voltage from 0v to 3v in 0.1v increments.

* set our plot scale (i.e. x axis to the n2 vector)
setscale n2 
* plotting properties
set title = 'DC Analysis: Current Output vs Drain Voltage' 
set xlabel = 'Drain Volage (V)'
set ylabel = 'Current Output (uA)'
set yhigh = 46
set ylow = 52
set filename = {$generic_prefix}{'_dc_analysis'}

gnuplot $filename (v2#branch*-1e+06) ylimit $ylow $yhigh title $title xlabel $xlabel ylabel $ylabel 

echo '* Writing all simulation data to a textfile'

set filetype=ascii
set filename = {$generic_prefix}{'_results.raw'}
write $filename

.ENDC
