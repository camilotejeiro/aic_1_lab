Four Transistor Current Mirror Simulation Testbench (DC)

* ---
* Netlist
* ---
.INCLUDE four_transistor_current_mirror_simulation_netlist.spice

* ---
* Control (Interactive Interpreter)
* ---
.CONTROL

    $ Make a directory for our output simulation files.
    shell mkdir -p results 
    $ Generic prefix for our output files
    set generic_prefix = 'results/four_transistor_current_mirror_simulation'
    
    $ Operating Point analysis $
    echo  '* Operating point analysis: Current match '

    OP                      
    print all               
    $ Output current over input current (with 1V load"): should be 1 for best match.
    print (v2#branch/v1#branch)

    $ DC Analysis
    $ ---
    echo '* DC analysis: Voltage dependence of current mirror'

    DC V2 0V 5V 0.1V          ; Sweep Collector voltage from 0v to 5V in 0.1v increments.

    $ Plotting
    $ ---
    $ plotting properties
    $ set our plot scale (i.e. x axis to the n2 vector)
    setscale n2 
    set title = 'DC Analysis: Current Output vs Collector Voltage' 
    set xlabel = 'Collector Volage (V)'
    set ylabel = 'Current Output (uA)'
    set yhigh = 51
    set ylow = 49
    set filename = {$generic_prefix}{'_analysis_dc'}
    gnuplot filename (v2#branch*-1e+06) ylimit $ylow $yhigh title $title xlabel $xlabel ylabel $ylabel 

    $ Write Simulation Data $
    echo '* Writing all simulation data to a textfile'

    set filetype=ascii
    set filename = {$generic_prefix}{'_results_dc.raw'}
    write $filename

.ENDC
