MOS Current Mirror With Cascode Stage Simulation Testbench (DC)

* ---
* Netlist
* ---
.INCLUDE mos_current_mirror_cascode_stage_simulation_netlist.spice

* ---
* Control (Interactive Interpreter)
* ---
.CONTROL

    $ Make a directory for our output simulation files.
    shell mkdir -p results 
    $ Generic prefix for our output files
    set generic_prefix = 'results/mos_current_mirror_cascode_stage_simulation'
    
    $ Operating Point analysis
    $ ---
    echo  '* Operating point analysis: Current match '

    OP                      
    print all               
    $ Output current over input current (with 1V load"): should be 1 for best match.
    print (v2#branch/v1#branch)

    $ DC Analysis
    $ ---
    echo '* DC analysis: Voltage dependence of current mirror'

    DC V2 0V 3V 0.1V          ; Sweep Drain voltage from 0v to 3V in 0.1v increments.

    $ Plotting
    $ ---
    $ plotting properties
    $ set our plot scale (i.e. x axis to the n2 vector)
    setscale n2 
    set title = 'DC Analysis: Current Output vs Drain Voltage' 
    set xlabel = 'Drain Voltage (V)'
    set ylabel = 'Current Output (uA)'
    set yhigh = 49.9
    set ylow = 49.1
    set filename = {$generic_prefix}{'_analysis_dc'}
    gnuplot $filename (v2#branch*-1e+06) ylimit $ylow $yhigh title $title xlabel $xlabel ylabel $ylabel 

    $ Write Simulation Data $
    echo '* Writing all simulation data to a textfile'

    set filetype=ascii
    set filename = {$generic_prefix}{'_results_dc.raw'}
    write $filename

.ENDC
