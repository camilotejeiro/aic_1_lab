* /media/camilo/data/workspaces/personal_projects/self_learning_courses/aic_1-analog_integrated_circuits/lab_assignments/2_simulation/ce_amplifier.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sun 20 Aug 2017 12:12:42 PM JST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
R4  /n2 /0 1KR		
R1  /n_pos /n1 100KR		
R2  /n1 /0 24KR		
R3  /n_pos /n_out 3.9KR		
C1  /n_in /n1 10uF		
V1  /n_pos /0 12V		
V2  /n_in /0 dc 0 ac 1.0 sin(0 1 1KHz)		
Q1  /n_out /n1 /n2 generic		;Node Sequence Spec.<c,b,e>

.end
