* /media/camilo/data/workspaces/academia/self_study/aic_1-analog_integrated_circuits/lab_assignments/3_current_mirrors/6_pnp_wilson_current_mirror/pnp_wilson_current_mirror.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Thu 21 Sep 2017 12:41:30 PM JST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
I1  /n3 /0 50uA		
V2  /n2 /0 4V		
V1  /n_pos /0 5V		
Q1  /n1 /n3 /n1 /n_pos PNP-Split-COLL		;Node Sequence Spec.<c1,c2,b,e>
Q2  /n2 /n3 /n1 PNP		;Node Sequence Spec.<c,b,e>

.end
