* Device Models

*      Name     Type(parameters) 
* ------------------------------
.MODEL generic  NPN

