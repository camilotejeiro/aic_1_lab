* Widely Used MOS Current Mirrors Simulation Netlist: 1st circuit (3-23) 
* Widely used mirror

* ---
* Subcircuits and Model parametters
* ---
.INCLUDE ../../device_parameter_libraries/cmos_hp_gmos10qa_350.spice
.INCLUDE ../../device_parameter_libraries/cmos_tsmc_cmos035_350.spice

* ---
* Netlist: Circuit Elements (Devices)
* ---
* dev <nets>            <values>
* -----------------------------------------------
V1    n_pos 0           3V		
I1    n_pos n3          50uA		
I2    n_pos n1          50uA	    
M1    n3    n3 0  0     hp_gmos10qa_n w=4u   l=2u   ; alternatively: tsmc_cmos_035n	
M2    n1    n3 n5 0     hp_gmos10qa_n w=100u l=2u 	
M3    n5    n1 0  0     hp_gmos10qa_n w=10u  l=5u 	
M4    n2    n3 n4 0     hp_gmos10qa_n w=100u l=2u 
M5    n4    n1 0  0     hp_gmos10qa_n w=10u  l=5u 
V2    n2    0           1V		

.END
