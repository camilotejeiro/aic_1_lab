* CMOS 0.350uM Process NMOS Devices Modified for Mismatch Monte-carlo Simulation

* ---
* Subcircuits and Model Parameters
* ---
* Note: we have included model declarations within each subcircuit to support 
* varying parameters for each transistor in the netlist individually 
* (for our missmatch Monte-carlo simulation).
* Otherwise: If we keep models "global" all parameter changes will be propagated 
* to all transistors in the netlist and the mismatch simulation won't work.

.SUBCKT hp_gmos10qa_n drain gate source bulk width=10u length=1u
* Nets: 1 (drain), 2 (gate), 3 (source), 4 (substrate/bulk)
* Values: Width and length of NMOS transistor.
* dev   <nets>                  model         <values>
* -----------------------------------------------------------
M1      drain gate source bulk  hp_gmos10qa_n w={width} l={length} 

.MODEL hp_gmos10qa_n NMOS ( level = 49 ; BSIM3 model 
+version = 3.3.0          tnom    = 27             tox     = 7.9e-9
+xj      = 1.5e-7         nch     = 1.7e17         vth0    = 0.5232192
+k1      = 0.6154629      k2      = 4.397909e-3    k3      = 49.5247378
+k3b     = 4.7261974      w0      = 1.428416e-5    nlx     = 1.990092e-7
+dvt0w   = 0              dvt1w   = 5.3e6          dvt2w   = -0.032
+dvt0    = 5.6285572      dvt1    = 0.8617134      dvt2    = -0.0569348
+u0      = 434.5143164    ua      = 1.066678e-10   ub      = 1.842089e-18
+uc      = 6.794094e-11   vsat    = 1.287889e5     a0      = 0.9907028
+ags     = 0.2642984      b0      = 1.894576e-6    b1      = 5e-6
+keta    = 1.06235e-3     a1      = 0              a2      = 1
+rdsw    = 976.0244735    prwg    = 2.031257e-3    prwb    = -1e-3
+wr      = 1              wint    = 5.506511e-8    lint    = 2.410167e-9
+xl      = -5e-8          xw      = 0              dwg     = -1.243637e-8
+dwb     = 5.537948e-9    voff    = -0.1310071     nfactor = 0.9944094
+cit     = 0              cdsc    = 1.527511e-3    cdscd   = 0
+cdscb   = 0              eta0    = 1.520266e-3    etab    = 0
+dsub    = 0.1067061      pclm    = 0.8764469      pdiblc1 = 0.5431391
+pdiblc2 = 4.15356e-3     pdiblcb = 0              drout   = 0.996452
+pscbe1  = 7.253118e9     pscbe2  = 5e-10          pvag    = 0.1772609
+delta   = 0.01           mobmod  = 1              prt     = 0
+ute     = -1.5           kt1     = -0.11          kt1l    = 0
+kt2     = 0.022          ua1     = 4.31e-9        ub1     = -7.61e-18
+uc1     = -5.6e-11       at      = 3.3e4          wl      = 0
+wln     = 1              ww      = 0              wwn     = 1
+wwl     = 0              ll      = 0              lln     = 1
+lw      = 0              lwn     = 1              lwl     = 0
+capmod  = 2              cgdo    = 3.97e-10       cgso    = 3.97e-10
+cgbo    = 0              cj      = 9.231271e-4    pb      = 0.8509074
+mj      = 0.3818435      cjsw    = 1.840483e-10   pbsw    = 0.9887463
+mjsw    = 0.1583859      pvth0   = -0.0115229     prdsw   = -139.443262
+pk2     = 3.497665e-4    wketa   = -1.09799e-3    lketa   = -7.09023e-3 )

.ENDS hp_gmos10qa_n

.SUBCKT tsmc_cmos_035n drain gate source bulk width=10u length=1u
* Nets: 1 (drain), 2 (gate), 3 (source), 4 (substrate/bulk)
* Values: Width and length of NMOS transistor.
* dev   <nets>                  model         <values>
* -----------------------------------------------------------
M1      drain gate source bulk  hp_gmos10qa_n w={width} l={length} 

.MODEL tsmc_cmos_035n NMOS ( level = 49 ; BSIM3 model 
+version = 3.3.0          tnom    = 27             tox     = 7.6e-9
+xj      = 1.5e-7         nch     = 1.7e17         vth0    = 0.4964448
+k1      = 0.5307769      k2      = 0.0199705      k3      = 0.2963637
+k3b     = 0.2012165      w0      = 2.836319e-6    nlx     = 2.894802e-7
+dvt0w   = 0              dvt1w   = 5.3e6          dvt2w   = -0.032
+dvt0    = 0.112017       dvt1    = 0.2453972      dvt2    = -0.171915
+u0      = 444.9381976    ua      = 2.921284e-10   ub      = 1.773281e-18
+uc      = 7.067896e-11   vsat    = 1.130785e5     a0      = 1.1356246
+ags     = 0.2810374      b0      = 2.844393e-7    b1      = 5e-6
+keta    = -7.8181e-3     a1      = 0              a2      = 1
+rdsw    = 925.2701982    prwg    = -1e-3          prwb    = -1e-3
+wr      = 1              wint    = 7.186965e-8    lint    = 1.735515e-9
+xl      = -2e-8          xw      = 0              dwg     = -1.712973e-8
+dwb     = 5.851691e-9    voff    = -0.132935      nfactor = 0.5710974
+cit     = 0              cdsc    = 8.607229e-4    cdscd   = 0
+cdscb   = 0              eta0    = 2.128321e-3    etab    = 0
+dsub    = 0.0257957      pclm    = 0.6766314      pdiblc1 = 1
+pdiblc2 = 1.787424e-3    pdiblcb = 0              drout   = 0.7873539
+pscbe1  = 6.973485e9     pscbe2  = 1.46235e-7     pvag    = 0.05
+delta   = 0.01           mobmod  = 1              prt     = 0
+ute     = -1.5           kt1     = -0.11          kt1l    = 0
+kt2     = 0.022          ua1     = 4.31e-9        ub1     = -7.61e-18
+uc1     = -5.6e-11       at      = 3.3e4          wl      = 0
+wln     = 1              ww      = 0              wwn     = 1
+wwl     = 0              ll      = 0              lln     = 1
+lw      = 0              lwn     = 1              lwl     = 0
+capmod  = 2              cgdo    = 1.96e-10       cgso    = 1.96e-10
+cgbo    = 0              cj      = 9.276962e-4    pb      = 0.8157962
+mj      = 0.3557696      cjsw    = 3.181055e-10   pbsw    = 0.6869149
+mjsw    = 0.1            pvth0   = -0.0252481     prdsw   = -96.4502805
+pk2     = -4.805372e-3   wketa   = -7.643187e-4   lketa   = -0.0129496 )

.ENDS tsmc_cmos_035n
