* Example from https://sourceforge.net/p/ngspice/discussion/133842/thread/5d3537b2/
* Taken as verbatim reference (untested)
* Thoroughly commented for understanding (feel free to remove comments).
* (exec-spice "ngspice -b %s" t)

* the model is within the subckt, so we have separate ones
* for each "inverter" instance

* ---
* Netlist: Circuit Elements (Devices)
* ---
* dev <nets>        <values>
* ------------------------------
vdd   vdd  0        DC=1.0
x1    out1 in1  vdd inverter
x2    out2 in2  vdd inverter
r1    in1  out1     2Meg
r2    in2  out2     2Meg

* ---
* Subcircuit and Included Models (for each created subcircuit instance)
* --- 
.SUBCKT inverter out in vdd
m1  out in  vdd vdd   pmos l=45n w=200n
m2  out in  0   0     nmos l=45n w=200n
.MODEL pmos pmos ( version=4.7 level=54 )
.MODEL nmos nmos ( version=4.7 level=54 )
.ENDS inverter

* ---
* Control block (interactive interpreter)
* ---
.CONTROL
define agauss(nom,avar,sig) (nom + avar/sig * sgauss(0))

OP

print v(out1) v(out2)

let vth0_x1 = agauss(0.8, 0.1, 3)
let vth0_x2 = agauss(0.8, 0.1, 3)

altermod x1:pmos vth0 vth0_x1
altermod x2:pmos vth0 vth0_x2

OP

print v(out1) v(out2)

showmod m.x1.m1 m.x2.m1

* you cant access a model parameter, only device parameters
*print @m.x1.m1[w]
*print @m.x1.m1[vth]


.ENDC
.END
