* /media/camilo/data/workspaces/academia/self_study/aic_1-analog_integrated_circuits/lab_assignments/3_current_mirrors/4_emitter_resistors_negative_feedback/emitter_resistors_negative_feedback.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Tue 19 Sep 2017 02:53:36 PM JST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: 
I1  n_pos n1 50uA		
Q1  n1 n1 n3 npn1		;Node Sequence Spec.<c,b,e>
Q2  n2 n1 n4 npn1		;Node Sequence Spec.<c,b,e>
V2  n2 0 1V		
V1  n_pos 0 5V		
R1  n3 0 6KR		
R2  n4 0 6KR		

.end
