Effecting a Monte Carlo calculation in ngspice
* Taken as verbatim reference from NGSPICE examples 
* Thoroughly commented for understanding (feel free to remove comments).

* ---
* Netlist
* ---
V1 N001 0 AC 1 DC 0
R1 N002 N001 141
 
C1 OUT 0 1e-09
L1 OUT 0 10e-06
C2 N002 0 1e-09
L2 N002 0 10e-06
L3 N003 N002 40e-06
C3 OUT N003 250e-12
 
R2 0 OUT 141

.CONTROL
    let mc_runs = 5
    let run = 0
    $ create a new plot
    set curplot=new          
    $ store its name to 'scratch'
    set scratch=$curplot     
    $ make 'scratch' the active plot 
    setplot $scratch         
    $ create a vector in plot 'scratch' to store bandwidth data
    let bwh=unitvec(mc_runs) 

    $ define distributions for random numbers:
    $ unif: uniform distribution, deviation relativ to nominal value
    $ aunif: uniform distribution, deviation absolut
    $ gauss: Gaussian distribution, deviation relativ to nominal value
    $ agauss: Gaussian distribution, deviation absolut
    $ limit: if unif. distributed value >=0 then add +avar to nom, else -avar
    define unif(nom, rvar) (nom + (nom*rvar) * sunif(0))
    define aunif(nom, avar) (nom + avar * sunif(0))
    define gauss(nom, rvar, sig) (nom + (nom*rvar)/sig * sgauss(0))
    define agauss(nom, avar, sig) (nom + avar/sig * sgauss(0))
    define limit(nom, avar) (nom + ((sgauss(0) >= 0) ? avar : -avar))

    dowhile run < mc_runs   
        alter c1 = unif(1e-09, 0.1)
        alter l1 = unif(10e-06, 0.1)
        alter c2 = unif(1e-09, 0.1)
        alter l2 = unif(10e-06, 0.1)
        alter l3 = unif(40e-06, 0.1)
        alter c3 = limit(250e-12, 25e-12)
         
        ac oct 100 250K 10Meg
         	
        $ measure bandwidth at -10 dB
        meas ac bw trig vdb(out) val=-10 rise=1 targ vdb(out) val=-10 fall=1
        $ create a variable from the vector  
        set run ="$&run"            
        $ store the current plot to dt
        set dt = $curplot           
        $ make 'scratch' the active plot
        setplot $scratch            
        $ store the output vector to plot 'scratch'
        let vout{$run}={$dt}.v(out) 
        $ store bw to vector bwh in plot 'scratch'
        let bwh[run]={$dt}.bw       
        $ go back to the previous plot
        setplot $dt                 
        let run = run + 1      	
    end   
       
    plot db({$scratch}.allv)
    echo
    print {$scratch}.bwh
.ENDC

.END
